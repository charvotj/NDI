library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity FDAC is
	
    Port ( CS_b : in  STD_LOGIC;
           SCLK : in  STD_LOGIC;
           fr_end : out  STD_LOGIC;
           fr_start : out  STD_LOGIC;
           fr_error : out  STD_LOGIC);
end FDAC;

architecture Behavioral of FDAC is

begin

    

end architecture;